# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__inv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  4.464000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.085000 1.550000 7.070000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.379200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.585000 1.920000 7.575000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.185000  0.085000 0.445000 1.130000 ;
      RECT 0.565000  1.330000 0.885000 2.995000 ;
      RECT 0.615000  0.350000 0.945000 1.130000 ;
      RECT 0.615000  1.130000 0.885000 1.330000 ;
      RECT 1.055000  1.940000 1.345000 3.245000 ;
      RECT 1.070000  1.350000 1.380000 1.770000 ;
      RECT 1.115000  0.085000 1.375000 1.130000 ;
      RECT 1.515000  1.940000 1.845000 2.980000 ;
      RECT 1.555000  0.350000 1.845000 1.940000 ;
      RECT 2.020000  1.350000 2.310000 1.770000 ;
      RECT 2.025000  0.085000 2.305000 1.130000 ;
      RECT 2.045000  1.940000 2.295000 3.245000 ;
      RECT 2.465000  1.940000 2.795000 2.980000 ;
      RECT 2.485000  0.350000 2.795000 1.940000 ;
      RECT 2.970000  1.350000 3.245000 1.770000 ;
      RECT 2.975000  0.085000 3.245000 1.130000 ;
      RECT 2.995000  1.940000 3.245000 3.245000 ;
      RECT 3.415000  0.350000 3.710000 2.980000 ;
      RECT 3.885000  1.350000 4.165000 1.770000 ;
      RECT 3.890000  0.085000 4.150000 1.130000 ;
      RECT 3.915000  1.940000 4.150000 3.245000 ;
      RECT 4.340000  0.350000 4.595000 1.940000 ;
      RECT 4.340000  1.940000 4.630000 2.980000 ;
      RECT 4.765000  0.085000 5.025000 1.130000 ;
      RECT 4.770000  1.350000 5.085000 1.770000 ;
      RECT 4.810000  1.940000 5.095000 3.245000 ;
      RECT 5.215000  0.350000 5.525000 1.180000 ;
      RECT 5.265000  1.180000 5.525000 1.285000 ;
      RECT 5.265000  1.285000 5.580000 2.980000 ;
      RECT 5.705000  0.085000 6.025000 1.130000 ;
      RECT 5.755000  1.350000 6.090000 1.770000 ;
      RECT 5.765000  1.940000 6.095000 3.245000 ;
      RECT 6.195000  0.350000 6.525000 1.180000 ;
      RECT 6.265000  1.180000 6.525000 1.285000 ;
      RECT 6.265000  1.285000 6.595000 2.980000 ;
      RECT 6.705000  0.085000 7.045000 1.130000 ;
      RECT 6.765000  1.940000 7.095000 3.245000 ;
      RECT 6.770000  1.350000 7.090000 1.770000 ;
      RECT 7.215000  0.350000 7.545000 1.130000 ;
      RECT 7.265000  1.130000 7.545000 2.980000 ;
      RECT 7.715000  0.085000 8.045000 1.130000 ;
      RECT 7.735000  1.820000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 0.645000  1.950000 0.815000 2.120000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.145000  1.580000 1.315000 1.750000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.950000 1.765000 2.120000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.085000  1.580000 2.255000 1.750000 ;
      RECT 2.545000  1.950000 2.715000 2.120000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.025000  1.580000 3.195000 1.750000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.495000  1.950000 3.665000 2.120000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.940000  1.580000 4.110000 1.750000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.395000  1.950000 4.565000 2.120000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.850000  1.580000 5.020000 1.750000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.345000  1.950000 5.515000 2.120000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.845000  1.580000 6.015000 1.750000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.345000  1.950000 6.515000 2.120000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.840000  1.580000 7.010000 1.750000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.345000  1.950000 7.515000 2.120000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ms__inv_16
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__or4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.470000 3.735000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.130000 4.395000 1.300000 ;
        RECT 2.525000 1.300000 3.235000 1.410000 ;
        RECT 2.615000 1.410000 3.235000 1.550000 ;
        RECT 4.065000 1.300000 4.395000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.605000 1.365000 6.285000 1.770000 ;
        RECT 4.925000 1.770000 6.285000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285000 0.255000 6.615000 0.855000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.326900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.945000 1.820000 ;
        RECT 0.125000 1.820000 2.275000 2.150000 ;
        RECT 0.615000 0.350000 0.945000 0.980000 ;
        RECT 0.615000 0.980000 1.945000 1.150000 ;
        RECT 0.615000 1.150000 0.945000 1.300000 ;
        RECT 0.615000 2.150000 0.845000 2.980000 ;
        RECT 1.515000 2.150000 1.745000 2.980000 ;
        RECT 1.615000 0.350000 1.945000 0.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  2.320000 0.445000 3.245000 ;
      RECT 1.015000  2.320000 1.345000 3.245000 ;
      RECT 1.115000  0.085000 1.445000 0.810000 ;
      RECT 1.315000  1.320000 2.325000 1.650000 ;
      RECT 1.915000  2.320000 2.245000 3.245000 ;
      RECT 2.155000  0.790000 5.100000 0.960000 ;
      RECT 2.155000  0.960000 2.325000 1.320000 ;
      RECT 2.380000  0.085000 2.740000 0.620000 ;
      RECT 2.475000  1.940000 2.805000 1.970000 ;
      RECT 2.475000  1.970000 4.675000 2.140000 ;
      RECT 2.475000  2.140000 2.805000 2.190000 ;
      RECT 2.475000  2.190000 2.755000 2.980000 ;
      RECT 2.920000  0.350000 3.250000 0.790000 ;
      RECT 2.925000  2.360000 4.175000 2.560000 ;
      RECT 2.925000  2.560000 3.205000 2.980000 ;
      RECT 3.375000  2.730000 3.705000 3.245000 ;
      RECT 3.430000  0.085000 4.590000 0.620000 ;
      RECT 3.825000  2.310000 4.175000 2.360000 ;
      RECT 3.895000  2.560000 4.175000 2.980000 ;
      RECT 4.345000  1.940000 4.675000 1.970000 ;
      RECT 4.345000  2.140000 4.675000 2.360000 ;
      RECT 4.345000  2.360000 6.575000 2.530000 ;
      RECT 4.345000  2.530000 4.675000 2.980000 ;
      RECT 4.770000  0.350000 5.100000 0.790000 ;
      RECT 4.770000  0.960000 5.100000 1.025000 ;
      RECT 4.770000  1.025000 6.635000 1.195000 ;
      RECT 4.845000  2.700000 6.075000 2.980000 ;
      RECT 5.270000  0.085000 6.115000 0.680000 ;
      RECT 5.295000  1.950000 6.635000 2.120000 ;
      RECT 5.295000  2.120000 5.625000 2.190000 ;
      RECT 6.245000  2.290000 6.575000 2.360000 ;
      RECT 6.245000  2.530000 6.575000 2.980000 ;
      RECT 6.465000  1.195000 6.635000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ms__or4_4
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__dlxtn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.270300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.265000 0.350000 6.615000 0.980000 ;
        RECT 6.265000 0.980000 8.035000 1.150000 ;
        RECT 6.315000 1.820000 8.035000 1.990000 ;
        RECT 6.315000 1.990000 6.645000 2.980000 ;
        RECT 7.295000 0.350000 7.545000 0.980000 ;
        RECT 7.315000 1.990000 8.035000 2.150000 ;
        RECT 7.315000 2.150000 7.545000 2.980000 ;
        RECT 7.805000 1.150000 8.035000 1.820000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.500000 1.315000 1.830000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.555000 0.445000 0.660000 ;
      RECT 0.115000  0.660000 1.315000 0.830000 ;
      RECT 0.115000  0.830000 0.795000 1.130000 ;
      RECT 0.135000  1.950000 0.795000 2.120000 ;
      RECT 0.135000  2.120000 0.465000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 0.490000 ;
      RECT 0.625000  1.130000 0.795000 1.950000 ;
      RECT 0.635000  2.290000 0.965000 3.245000 ;
      RECT 1.135000  1.000000 1.885000 1.330000 ;
      RECT 1.135000  2.100000 1.655000 2.390000 ;
      RECT 1.135000  2.390000 3.160000 2.560000 ;
      RECT 1.135000  2.560000 1.655000 2.980000 ;
      RECT 1.145000  0.255000 2.645000 0.425000 ;
      RECT 1.145000  0.425000 1.315000 0.660000 ;
      RECT 1.485000  0.760000 1.885000 1.000000 ;
      RECT 1.485000  1.330000 1.885000 1.770000 ;
      RECT 1.485000  1.770000 1.655000 2.100000 ;
      RECT 1.825000  1.940000 2.225000 2.220000 ;
      RECT 2.055000  0.595000 2.305000 1.720000 ;
      RECT 2.055000  1.720000 3.540000 1.890000 ;
      RECT 2.055000  1.890000 2.225000 1.940000 ;
      RECT 2.360000  2.730000 2.820000 3.245000 ;
      RECT 2.475000  0.425000 2.645000 1.220000 ;
      RECT 2.475000  1.220000 3.000000 1.550000 ;
      RECT 2.815000  0.085000 3.145000 1.050000 ;
      RECT 2.990000  2.560000 3.160000 2.905000 ;
      RECT 2.990000  2.905000 4.220000 3.075000 ;
      RECT 3.210000  1.470000 3.540000 1.720000 ;
      RECT 3.315000  0.255000 4.445000 0.505000 ;
      RECT 3.315000  0.505000 3.485000 1.470000 ;
      RECT 3.360000  2.060000 3.880000 2.735000 ;
      RECT 3.655000  0.725000 4.720000 1.055000 ;
      RECT 3.710000  1.055000 3.880000 2.060000 ;
      RECT 4.050000  1.405000 4.380000 1.735000 ;
      RECT 4.050000  1.735000 4.220000 2.905000 ;
      RECT 4.390000  1.975000 5.830000 1.990000 ;
      RECT 4.390000  1.990000 5.645000 2.305000 ;
      RECT 4.390000  2.590000 5.145000 3.245000 ;
      RECT 4.550000  1.055000 4.720000 1.320000 ;
      RECT 4.550000  1.320000 5.490000 1.650000 ;
      RECT 4.890000  0.085000 5.140000 1.055000 ;
      RECT 5.315000  1.820000 5.830000 1.975000 ;
      RECT 5.315000  2.305000 5.645000 2.980000 ;
      RECT 5.320000  0.375000 5.570000 0.980000 ;
      RECT 5.320000  0.980000 5.830000 1.150000 ;
      RECT 5.660000  1.150000 5.830000 1.320000 ;
      RECT 5.660000  1.320000 7.490000 1.650000 ;
      RECT 5.660000  1.650000 5.830000 1.820000 ;
      RECT 5.750000  0.085000 6.080000 0.810000 ;
      RECT 5.815000  2.160000 6.145000 3.245000 ;
      RECT 6.785000  0.085000 7.115000 0.810000 ;
      RECT 6.815000  2.160000 7.145000 3.245000 ;
      RECT 7.715000  0.085000 8.045000 0.810000 ;
      RECT 7.715000  2.320000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ms__dlxtn_4
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__dfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725000 2.050000 2.055000 2.380000 ;
        RECT 1.885000 1.150000 2.275000 1.480000 ;
        RECT 1.885000 1.480000 2.055000 2.050000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.745000 2.030000 8.105000 2.980000 ;
        RECT 7.765000 0.350000 8.105000 1.130000 ;
        RECT 7.935000 1.130000 8.105000 2.030000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 1.135000 1.130000 ;
      RECT 0.115000  1.950000 0.845000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.545000  0.085000 0.795000 0.790000 ;
      RECT 0.645000  2.290000 0.815000 3.245000 ;
      RECT 0.675000  1.130000 1.135000 1.550000 ;
      RECT 0.675000  1.550000 0.845000 1.950000 ;
      RECT 0.965000  0.255000 1.815000 0.425000 ;
      RECT 0.965000  0.425000 1.135000 0.960000 ;
      RECT 1.015000  1.720000 1.475000 2.625000 ;
      RECT 1.015000  2.625000 2.275000 2.755000 ;
      RECT 1.015000  2.755000 4.990000 2.795000 ;
      RECT 1.015000  2.795000 1.345000 2.980000 ;
      RECT 1.305000  0.595000 1.475000 1.350000 ;
      RECT 1.305000  1.350000 1.715000 1.720000 ;
      RECT 1.575000  2.965000 1.935000 3.245000 ;
      RECT 1.645000  0.425000 1.815000 0.810000 ;
      RECT 1.645000  0.810000 2.520000 0.980000 ;
      RECT 1.985000  0.085000 2.180000 0.640000 ;
      RECT 2.105000  2.795000 3.540000 2.925000 ;
      RECT 2.225000  1.650000 2.615000 1.820000 ;
      RECT 2.225000  1.820000 2.555000 2.455000 ;
      RECT 2.350000  0.255000 3.755000 0.425000 ;
      RECT 2.350000  0.425000 2.520000 0.810000 ;
      RECT 2.445000  1.150000 2.860000 1.320000 ;
      RECT 2.445000  1.320000 2.615000 1.650000 ;
      RECT 2.690000  0.595000 2.860000 1.150000 ;
      RECT 2.755000  2.125000 2.955000 2.255000 ;
      RECT 2.755000  2.255000 4.135000 2.425000 ;
      RECT 2.755000  2.425000 2.955000 2.585000 ;
      RECT 2.785000  1.490000 3.200000 1.660000 ;
      RECT 2.785000  1.660000 2.955000 2.125000 ;
      RECT 3.030000  0.615000 3.415000 0.945000 ;
      RECT 3.030000  0.945000 3.200000 1.490000 ;
      RECT 3.140000  1.830000 3.540000 2.085000 ;
      RECT 3.370000  1.285000 3.755000 1.455000 ;
      RECT 3.370000  1.455000 3.540000 1.830000 ;
      RECT 3.370000  2.625000 4.990000 2.755000 ;
      RECT 3.585000  0.425000 3.755000 0.690000 ;
      RECT 3.585000  0.690000 4.575000 0.860000 ;
      RECT 3.585000  0.860000 3.755000 1.285000 ;
      RECT 3.710000  2.965000 4.100000 3.245000 ;
      RECT 3.925000  1.030000 4.915000 1.200000 ;
      RECT 3.925000  1.200000 4.650000 1.415000 ;
      RECT 3.965000  1.625000 4.310000 1.955000 ;
      RECT 3.965000  1.955000 4.135000 2.255000 ;
      RECT 3.985000  0.085000 4.235000 0.520000 ;
      RECT 4.305000  2.125000 4.650000 2.455000 ;
      RECT 4.405000  0.255000 5.890000 0.425000 ;
      RECT 4.405000  0.425000 4.575000 0.690000 ;
      RECT 4.480000  1.415000 4.650000 2.125000 ;
      RECT 4.745000  0.595000 5.075000 0.945000 ;
      RECT 4.745000  0.945000 4.915000 1.030000 ;
      RECT 4.820000  1.370000 5.415000 1.540000 ;
      RECT 4.820000  1.540000 4.990000 2.625000 ;
      RECT 4.820000  2.795000 4.990000 2.905000 ;
      RECT 4.820000  2.905000 5.875000 3.075000 ;
      RECT 5.085000  1.150000 5.415000 1.370000 ;
      RECT 5.160000  1.710000 5.755000 1.880000 ;
      RECT 5.160000  1.880000 5.330000 2.735000 ;
      RECT 5.245000  0.695000 5.755000 0.945000 ;
      RECT 5.545000  2.050000 5.875000 2.905000 ;
      RECT 5.560000  0.425000 5.890000 0.510000 ;
      RECT 5.585000  0.945000 5.755000 1.230000 ;
      RECT 5.585000  1.230000 7.240000 1.400000 ;
      RECT 5.585000  1.400000 5.755000 1.710000 ;
      RECT 6.085000  1.570000 6.415000 1.690000 ;
      RECT 6.085000  1.690000 7.765000 1.860000 ;
      RECT 6.085000  1.860000 6.415000 2.240000 ;
      RECT 6.225000  0.085000 6.555000 1.060000 ;
      RECT 6.235000  2.520000 6.565000 3.245000 ;
      RECT 6.785000  0.350000 7.115000 0.850000 ;
      RECT 6.785000  0.850000 7.595000 1.020000 ;
      RECT 6.790000  1.860000 7.040000 2.860000 ;
      RECT 6.910000  1.190000 7.240000 1.230000 ;
      RECT 6.910000  1.400000 7.240000 1.520000 ;
      RECT 7.240000  2.030000 7.570000 3.245000 ;
      RECT 7.300000  0.085000 7.595000 0.680000 ;
      RECT 7.425000  1.020000 7.595000 1.350000 ;
      RECT 7.425000  1.350000 7.765000 1.690000 ;
      RECT 8.275000  0.085000 8.525000 1.130000 ;
      RECT 8.275000  1.820000 8.525000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ms__dfxtp_2
END LIBRARY

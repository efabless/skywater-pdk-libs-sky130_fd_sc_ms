# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a221o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 1.450000 2.275000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.365000 1.260000 1.765000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 1.450000 2.760000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.180000 3.695000 1.550000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 1.180000 4.195000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.960000 0.855000 1.130000 ;
        RECT 0.100000 1.130000 0.335000 1.800000 ;
        RECT 0.100000 1.800000 0.930000 1.970000 ;
        RECT 0.600000 1.970000 0.930000 2.980000 ;
        RECT 0.605000 0.350000 0.855000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.150000  2.140000 0.400000 3.245000 ;
      RECT 0.175000  0.085000 0.425000 0.790000 ;
      RECT 0.525000  1.300000 1.195000 1.630000 ;
      RECT 1.025000  0.920000 4.220000 1.010000 ;
      RECT 1.025000  1.010000 3.100000 1.090000 ;
      RECT 1.025000  1.090000 1.195000 1.300000 ;
      RECT 1.035000  0.085000 1.560000 0.750000 ;
      RECT 1.130000  1.950000 1.380000 3.245000 ;
      RECT 1.565000  1.950000 2.730000 2.060000 ;
      RECT 1.565000  2.060000 3.315000 2.120000 ;
      RECT 1.565000  2.120000 1.815000 2.980000 ;
      RECT 2.015000  2.290000 2.345000 3.245000 ;
      RECT 2.020000  0.350000 2.890000 0.840000 ;
      RECT 2.020000  0.840000 4.220000 0.920000 ;
      RECT 2.020000  1.090000 3.100000 1.130000 ;
      RECT 2.535000  2.400000 2.785000 2.905000 ;
      RECT 2.535000  2.905000 3.685000 3.075000 ;
      RECT 2.540000  2.120000 3.315000 2.230000 ;
      RECT 2.930000  1.130000 3.100000 1.720000 ;
      RECT 2.930000  1.720000 4.215000 1.890000 ;
      RECT 2.985000  2.230000 3.315000 2.735000 ;
      RECT 3.350000  0.085000 3.720000 0.670000 ;
      RECT 3.515000  2.060000 3.685000 2.905000 ;
      RECT 3.885000  1.890000 4.215000 2.980000 ;
      RECT 3.890000  0.350000 4.220000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__a221o_2
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__mux2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 1.195000 1.550000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.470000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.450000 2.385000 1.780000 ;
        RECT 2.215000 1.130000 3.455000 1.300000 ;
        RECT 2.215000 1.300000 2.385000 1.450000 ;
        RECT 3.125000 1.300000 3.455000 1.460000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 0.770000 4.665000 2.140000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  1.825000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.905000 3.075000 ;
      RECT 0.170000  0.290000 2.750000 0.460000 ;
      RECT 0.170000  0.460000 0.500000 1.010000 ;
      RECT 0.620000  1.820000 1.535000 1.970000 ;
      RECT 0.620000  1.970000 3.165000 2.140000 ;
      RECT 0.620000  2.140000 0.840000 2.725000 ;
      RECT 0.670000  0.680000 1.535000 1.010000 ;
      RECT 1.015000  2.310000 2.825000 2.480000 ;
      RECT 1.015000  2.480000 1.345000 2.735000 ;
      RECT 1.365000  1.010000 1.535000 1.820000 ;
      RECT 1.575000  2.650000 1.905000 2.905000 ;
      RECT 1.715000  0.790000 3.170000 0.960000 ;
      RECT 1.715000  0.960000 2.045000 1.130000 ;
      RECT 2.075000  2.650000 2.405000 3.245000 ;
      RECT 2.420000  0.460000 2.750000 0.620000 ;
      RECT 2.555000  1.470000 2.885000 1.630000 ;
      RECT 2.555000  1.630000 3.795000 1.800000 ;
      RECT 2.575000  2.480000 2.825000 2.980000 ;
      RECT 2.995000  2.140000 3.165000 2.310000 ;
      RECT 2.995000  2.310000 5.165000 2.480000 ;
      RECT 3.000000  0.085000 3.170000 0.790000 ;
      RECT 3.335000  1.800000 3.795000 2.140000 ;
      RECT 3.340000  0.350000 3.670000 0.770000 ;
      RECT 3.340000  0.770000 3.795000 0.940000 ;
      RECT 3.625000  0.940000 3.795000 1.630000 ;
      RECT 3.840000  0.085000 4.230000 0.600000 ;
      RECT 3.870000  2.650000 4.210000 3.245000 ;
      RECT 4.780000  2.650000 5.165000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 1.130000 ;
      RECT 4.835000  1.300000 5.165000 2.310000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_ms__mux2_2
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a21bo_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.655000 1.450000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 0.435000 0.670000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.180000 2.845000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295000 0.350000 3.755000 1.130000 ;
        RECT 3.430000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.130000  1.940000 0.460000 1.950000 ;
      RECT 0.130000  1.950000 1.390000 2.120000 ;
      RECT 0.130000  2.120000 0.460000 2.980000 ;
      RECT 0.155000  0.840000 0.775000 1.095000 ;
      RECT 0.155000  1.095000 0.485000 1.340000 ;
      RECT 0.605000  0.085000 0.775000 0.840000 ;
      RECT 0.660000  2.290000 0.860000 3.245000 ;
      RECT 0.945000  0.660000 1.315000 1.110000 ;
      RECT 0.945000  1.110000 1.745000 1.280000 ;
      RECT 1.060000  2.120000 1.390000 2.980000 ;
      RECT 1.485000  0.085000 1.815000 0.930000 ;
      RECT 1.575000  1.280000 1.745000 1.940000 ;
      RECT 1.575000  1.940000 1.760000 2.240000 ;
      RECT 1.575000  2.240000 3.255000 2.410000 ;
      RECT 1.575000  2.410000 1.760000 2.980000 ;
      RECT 1.915000  1.100000 2.245000 1.770000 ;
      RECT 2.075000  0.350000 2.720000 0.940000 ;
      RECT 2.075000  0.940000 2.245000 1.100000 ;
      RECT 2.075000  1.770000 2.245000 1.820000 ;
      RECT 2.075000  1.820000 2.695000 2.070000 ;
      RECT 2.900000  0.085000 3.115000 0.895000 ;
      RECT 2.900000  2.580000 3.230000 3.245000 ;
      RECT 3.085000  1.320000 3.415000 1.650000 ;
      RECT 3.085000  1.650000 3.255000 2.240000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_ms__a21bo_1
END LIBRARY
